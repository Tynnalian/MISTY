//---------------------------------------------------------
// Class: axis_misty_params_pkg
//---------------------------------------------------------

// AXI-Stream ALU verification package.

package axis_misty_params_pkg;

    // Import UVM package.


parameter WIDTH = 200;


endpackage