//---------------------------------------------------------
// Interface: reset_intf
//---------------------------------------------------------

// Reset interface

interface reset_intf (
    input logic clk_i
);

    // Interface wires

    logic reset;

endinterface
