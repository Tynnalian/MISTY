//---------------------------------------------------------
// Class: MISTY_dv_pkg
//---------------------------------------------------------

// Verification package

package misty_pkg; 
   
    import pysv::*;
    import uvm_pkg::*;
    `include "uvm_macros.svh" 
    
    `include "misty_seq_item.sv"
    `include "misty_driver.sv"
    `include "misty_monitor.sv"
    `include "misty_agent.sv"
    `include "misty_cov.sv"
    `include "misty_scoreboard.sv"
endpackage