//---------------------------------------------------------
// Class: misty_top_pkg
//---------------------------------------------------------

// misty top verification package.

package misty_top_pkg;


    import uvm_pkg::*;
    import pysv::*;
    import misty_pkg::*;
    import reset_agent_pkg::*;
    
    parameter DURATION = 293;

    `include "uvm_macros.svh"
    `include "misty_seq_lib.sv"
    `include "misty_top_scoreboard.sv"
    `include "misty_env.sv"
    `include "misty_test.sv"

endpackage